library ieee;
use ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

entity instrMemory is port (
    Addr : in std_logic_vector(3 downto 0);
    C : out std_logic_vector(31 downto 0));
end instrMemory;

architecture arch1 of instrMemory is
    type instr_array is array (0 to 15) of std_logic_vector (31 downto 0);
    constant instrmem: instr_array := (
    "11111111111111111111111111111111", -- 0
    "10001010100101010101000011101111", -- 1
    "11111111111111111111111111111111", -- 2
    "00000000000000000000000000000000", -- 3
    "11111111111111111111111111111111", -- 4
    "00000000000000000000000000000000", -- 5
    "00000000101001100010000000100000", -- 6
    "11111111111111111111111111111111", -- 7
    "11111111111111111111111111111111", -- 8
    "11111111111111111111111111111111", -- 9
    "10101010101011110000101110001010", --10
    "11111111111111100000000000000000", --11
    "10001011101010111010111101010111", --12
    "11111111111111111111111111111111", --13
    "10110111000111010101010101111111", --14
    "11111111111111111111111111111111");--15
begin
    C <= instrmem(to_integer(unsigned(Addr)));
end arch1;